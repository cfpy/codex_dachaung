//�򵥵��ۼ�ģ��
`timescale 1ns/1ps
module read_write(
input clk,//ʱ��
input rst,//��λ
input [4:0]add1,//����ļ���

output reg [4:0]sum//������ܺ�
);
initial sum=5'h0;
always@(posedge clk,negedge rst)
begin
	if(!rst)
		begin
			sum<=5'h0;	
		end
	else
		begin
			sum<=sum + add1;
		end
end
endmodule 